library ieee;
use ieee.std_logic_1164.all;

entity praktiskt_prov_tb is
end entity;

architecture tb of praktiskt_prov_tb is

signal clk_s : std_logic;

begin
end;